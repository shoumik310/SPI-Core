module SPI ();

endmodule